module RVArch(
  input   clock,
  input   reset
);
endmodule
